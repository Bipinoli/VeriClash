module CircularStack ();

endmodule